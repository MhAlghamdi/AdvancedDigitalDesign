`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:29:32 02/27/2017 
// Design Name: 
// Module Name:    counter 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module counter(
    input wire clk, reset,
    input wire inc, dec,
    output reg [7:0] occupancy
    );
	
	
	reg [7:0] count = 0;
	
	always@(posedge clk) begin
		if (reset)
			count <= 0;
		else if (inc)
			count <= count + 1;
		else if (dec)
			count <= count - 1;
	end
	
	always @(*) begin
		occupancy = count;
	end
	
endmodule
